interface mem_intfc;
    bit start,write;
    logic [2:0] 