interface counter_if(input bit clk );
bit  rst ;
logic [3:0]count;

endinterface