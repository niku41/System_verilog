`timescale 1ns / 1ps
interface melay_0101_if();
bit rst;
bit clk;
logic seq_in;
logic seq_out;
endinterface